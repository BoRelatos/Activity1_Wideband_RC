* Wideband RC Voltage Divider
.options savecurrents

* Main Circuit
R1 in out 8.2e+06
R2 out 0 180000
C1 in out 0.0856p
C2 out 0 3.900p

* Variations
R1a in outa 8.2e+06
R2a outa 0 180000
C1a in outa 0.07704p
C2a outa 0 3.900p

R1b in outb 8.2e+06
R2b outb 0 180000
C1b in outb 0.09416p
C2b outb 0 3.900p

V1 in 0 pulse(-0.1 0.1 0 0.1u 0.1u 5u 10u) dc 1 ac 1

.control
  ac dec 10 1 1G
  wrdata output_ac.dat v(out) v(outa) v(outb)
  
  tran 0.01u 30u
  wrdata output_tran.dat v(out) v(outa) v(outb)
  quit
.endc
.end
